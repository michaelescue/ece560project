bind darkriscv darkriscv_checker_sva mychecker(CLK, RES, HLT, IDATA, DATAI);

